module test_multiplier;

endmodule
module test_multiplier

